-- megafunction wizard: %SRAM/SSRAM Controller v13.0%
-- GENERATION: XML
-- sramController.vhd

-- Generated using ACDS version 13.0sp1 232 at 2020.01.22.17:22:24

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sramController is
	port (
		clk           : in    std_logic                     := '0';             --        clock_reset.clk
		reset         : in    std_logic                     := '0';             --  clock_reset_reset.reset
		SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => '0'); -- external_interface.export
		SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    --                   .export
		SRAM_LB_N     : out   std_logic;                                        --                   .export
		SRAM_UB_N     : out   std_logic;                                        --                   .export
		SRAM_CE_N     : out   std_logic;                                        --                   .export
		SRAM_OE_N     : out   std_logic;                                        --                   .export
		SRAM_WE_N     : out   std_logic;                                        --                   .export
		address       : in    std_logic_vector(19 downto 0) := (others => '0'); --  avalon_sram_slave.address
		byteenable    : in    std_logic_vector(1 downto 0)  := (others => '0'); --                   .byteenable
		read          : in    std_logic                     := '0';             --                   .read
		write         : in    std_logic                     := '0';             --                   .write
		writedata     : in    std_logic_vector(15 downto 0) := (others => '0'); --                   .writedata
		readdata      : out   std_logic_vector(15 downto 0);                    --                   .readdata
		readdatavalid : out   std_logic                                         --                   .readdatavalid
	);
end entity sramController;

architecture rtl of sramController is
	component sramController_0002 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(31 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(31 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component sramController_0002;

begin

	sramcontroller_inst : component sramController_0002
		port map (
			clk           => clk,           --        clock_reset.clk
			reset         => reset,         --  clock_reset_reset.reset
			SRAM_DQ       => SRAM_DQ,       -- external_interface.export
			SRAM_ADDR     => SRAM_ADDR,     --                   .export
			SRAM_LB_N     => SRAM_LB_N,     --                   .export
			SRAM_UB_N     => SRAM_UB_N,     --                   .export
			SRAM_CE_N     => SRAM_CE_N,     --                   .export
			SRAM_OE_N     => SRAM_OE_N,     --                   .export
			SRAM_WE_N     => SRAM_WE_N,     --                   .export
			address       => address,       --  avalon_sram_slave.address
			byteenable    => byteenable,    --                   .byteenable
			read          => read,          --                   .read
			write         => write,         --                   .write
			writedata     => writedata,     --                   .writedata
			readdata      => readdata,      --                   .readdata
			readdatavalid => readdatavalid  --                   .readdatavalid
		);

end architecture rtl; -- of sramController
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2020 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_up_avalon_sram" version="13.0" >
-- Retrieval info: 	<generic name="board" value="DE2-115" />
-- Retrieval info: 	<generic name="pixel_buffer" value="false" />
-- Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
-- Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone IV E" />
-- Retrieval info: </instance>
-- IPFS_FILES : sramController.vho
-- RELATED_FILES: sramController.vhd, sramController_0002.v
